 `timescale 1ns/1ns
module BarrelShifter16bit(input [15:0] a ,input[3:0] s,output [15:0] sh );
   MUX16to1 MUX1 (.J({a[15],a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14]}),.s(s),.w(sh[15])),
            MUX2 (.J({a[14],a[15],a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13]}),.s(s),.w(sh[14])), 
            MUX3 (.J({a[13],a[14],a[15],a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12]}),.s(s),.w(sh[13])),
            MUX4 (.J({a[12],a[13],a[14],a[15],a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11]}),.s(s),.w(sh[12])),
            MUX5 (.J({a[11],a[12],a[13],a[14],a[15],a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10]}),.s(s),.w(sh[11])),
            MUX6 (.J({a[10],a[11],a[12],a[13],a[14],a[15],a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9]}),.s(s),.w(sh[10])),
            MUX7 (.J({a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8]}),.s(s),.w(sh[9])),
            MUX8 (.J({a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7]}),.s(s),.w(sh[8])),
            MUX9 (.J({a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[0],a[1],a[2],a[3],a[4],a[5],a[6]}),.s(s),.w(sh[7])),
            MUX10 (.J({a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[0],a[1],a[2],a[3],a[4],a[5]}),.s(s),.w(sh[6])),
            MUX11 (.J({a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[0],a[1],a[2],a[3],a[4]}),.s(s),.w(sh[5])),
            MUX12 (.J({a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[0],a[1],a[2],a[3]}),.s(s),.w(sh[4])),
            MUX13 (.J({a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[0],a[1],a[2]}),.s(s),.w(sh[3])),
            MUX14 (.J({a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[0],a[1]}),.s(s),.w(sh[2])),
            MUX15 (.J({a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15],a[0]}),.s(s),.w(sh[1])),
            MUX16 (.J({a[0],a[1],a[2],a[3],a[4],a[5],a[6],a[7],a[8],a[9],a[10],a[11],a[12],a[13],a[14],a[15]}),.s(s),.w(sh[0]));
endmodule